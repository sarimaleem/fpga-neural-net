`ifndef GLOBAL_PARAMS_VH
`define GLOBAL_PARAMS_VH

parameter HEIGHT = 20;
parameter LENGTH = 30;

`endif