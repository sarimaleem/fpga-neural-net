`ifndef GLOBAL_PARAMS_VH
`define GLOBAL_PARAMS_VH

parameter WIDTH = 200;
parameter HEIGHT = 300;

`endif