`ifndef GLOBAL_PARAMS_VH
`define GLOBAL_PARAMS_VH

parameter LENGTH = 20;
parameter WIDTH = 30;

parameter SHIFT = LENGTH / 10;
parameter LEFT = LENGTH * 4 / 10;

parameter LOWER_GREEN_ONE = 18;
parameter LOWER_GREEN_TWO = 25;
parameter LOWER_GREEN_THREE = 25;

parameter UPPER_GREEN_ONE = 43;
parameter UPPER_GREEN_TWO = 255;
parameter UPPER_GREEN_THREE = 255;

`endif