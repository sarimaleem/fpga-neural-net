module data_init (inout logic [7:0] image [{LENGTH-1}:0][{WIDTH-1}:0]);

logic [7:0] image [19:0][29:0];

initial begin
    image[0][0][0] = 8'd40;
    image[0][0][1] = 8'd122;
    image[0][0][2] = 8'd34;
    image[0][1][0] = 8'd40;
    image[0][1][1] = 8'd123;
    image[0][1][2] = 8'd33;
    image[0][2][0] = 8'd42;
    image[0][2][1] = 8'd125;
    image[0][2][2] = 8'd34;
    image[0][3][0] = 8'd45;
    image[0][3][1] = 8'd130;
    image[0][3][2] = 8'd37;
    image[0][4][0] = 8'd45;
    image[0][4][1] = 8'd130;
    image[0][4][2] = 8'd37;
    image[0][5][0] = 8'd45;
    image[0][5][1] = 8'd132;
    image[0][5][2] = 8'd36;
    image[0][6][0] = 8'd48;
    image[0][6][1] = 8'd135;
    image[0][6][2] = 8'd38;
    image[0][7][0] = 8'd49;
    image[0][7][1] = 8'd137;
    image[0][7][2] = 8'd39;
    image[0][8][0] = 8'd50;
    image[0][8][1] = 8'd139;
    image[0][8][2] = 8'd42;
    image[0][9][0] = 8'd51;
    image[0][9][1] = 8'd141;
    image[0][9][2] = 8'd40;
    image[0][10][0] = 8'd52;
    image[0][10][1] = 8'd143;
    image[0][10][2] = 8'd41;
    image[0][11][0] = 8'd52;
    image[0][11][1] = 8'd143;
    image[0][11][2] = 8'd42;
    image[0][12][0] = 8'd54;
    image[0][12][1] = 8'd144;
    image[0][12][2] = 8'd42;
    image[0][13][0] = 8'd53;
    image[0][13][1] = 8'd144;
    image[0][13][2] = 8'd42;
    image[0][14][0] = 8'd52;
    image[0][14][1] = 8'd144;
    image[0][14][2] = 8'd42;
    image[0][15][0] = 8'd53;
    image[0][15][1] = 8'd145;
    image[0][15][2] = 8'd43;
    image[0][16][0] = 8'd53;
    image[0][16][1] = 8'd144;
    image[0][16][2] = 8'd43;
    image[0][17][0] = 8'd53;
    image[0][17][1] = 8'd145;
    image[0][17][2] = 8'd44;
    image[0][18][0] = 8'd54;
    image[0][18][1] = 8'd145;
    image[0][18][2] = 8'd45;
    image[0][19][0] = 8'd53;
    image[0][19][1] = 8'd142;
    image[0][19][2] = 8'd43;
    image[0][20][0] = 8'd51;
    image[0][20][1] = 8'd141;
    image[0][20][2] = 8'd42;
    image[0][21][0] = 8'd51;
    image[0][21][1] = 8'd140;
    image[0][21][2] = 8'd42;
    image[0][22][0] = 8'd49;
    image[0][22][1] = 8'd138;
    image[0][22][2] = 8'd41;
    image[0][23][0] = 8'd48;
    image[0][23][1] = 8'd136;
    image[0][23][2] = 8'd41;
    image[0][24][0] = 8'd47;
    image[0][24][1] = 8'd135;
    image[0][24][2] = 8'd41;
    image[0][25][0] = 8'd47;
    image[0][25][1] = 8'd135;
    image[0][25][2] = 8'd42;
    image[0][26][0] = 8'd42;
    image[0][26][1] = 8'd130;
    image[0][26][2] = 8'd41;
    image[0][27][0] = 8'd42;
    image[0][27][1] = 8'd128;
    image[0][27][2] = 8'd38;
    image[0][28][0] = 8'd40;
    image[0][28][1] = 8'd126;
    image[0][28][2] = 8'd39;
    image[0][29][0] = 8'd39;
    image[0][29][1] = 8'd123;
    image[0][29][2] = 8'd37;
    image[1][0][0] = 8'd43;
    image[1][0][1] = 8'd127;
    image[1][0][2] = 8'd32;
    image[1][1][0] = 8'd41;
    image[1][1][1] = 8'd127;
    image[1][1][2] = 8'd31;
    image[1][2][0] = 8'd45;
    image[1][2][1] = 8'd131;
    image[1][2][2] = 8'd33;
    image[1][3][0] = 8'd43;
    image[1][3][1] = 8'd132;
    image[1][3][2] = 8'd33;
    image[1][4][0] = 8'd47;
    image[1][4][1] = 8'd135;
    image[1][4][2] = 8'd34;
    image[1][5][0] = 8'd49;
    image[1][5][1] = 8'd138;
    image[1][5][2] = 8'd35;
    image[1][6][0] = 8'd51;
    image[1][6][1] = 8'd141;
    image[1][6][2] = 8'd37;
    image[1][7][0] = 8'd51;
    image[1][7][1] = 8'd141;
    image[1][7][2] = 8'd36;
    image[1][8][0] = 8'd51;
    image[1][8][1] = 8'd143;
    image[1][8][2] = 8'd38;
    image[1][9][0] = 8'd52;
    image[1][9][1] = 8'd144;
    image[1][9][2] = 8'd36;
    image[1][10][0] = 8'd53;
    image[1][10][1] = 8'd147;
    image[1][10][2] = 8'd39;
    image[1][11][0] = 8'd52;
    image[1][11][1] = 8'd146;
    image[1][11][2] = 8'd38;
    image[1][12][0] = 8'd53;
    image[1][12][1] = 8'd147;
    image[1][12][2] = 8'd39;
    image[1][13][0] = 8'd52;
    image[1][13][1] = 8'd147;
    image[1][13][2] = 8'd38;
    image[1][14][0] = 8'd52;
    image[1][14][1] = 8'd147;
    image[1][14][2] = 8'd39;
    image[1][15][0] = 8'd54;
    image[1][15][1] = 8'd150;
    image[1][15][2] = 8'd41;
    image[1][16][0] = 8'd56;
    image[1][16][1] = 8'd149;
    image[1][16][2] = 8'd41;
    image[1][17][0] = 8'd55;
    image[1][17][1] = 8'd148;
    image[1][17][2] = 8'd43;
    image[1][18][0] = 8'd55;
    image[1][18][1] = 8'd148;
    image[1][18][2] = 8'd43;
    image[1][19][0] = 8'd55;
    image[1][19][1] = 8'd146;
    image[1][19][2] = 8'd43;
    image[1][20][0] = 8'd53;
    image[1][20][1] = 8'd144;
    image[1][20][2] = 8'd41;
    image[1][21][0] = 8'd51;
    image[1][21][1] = 8'd142;
    image[1][21][2] = 8'd40;
    image[1][22][0] = 8'd53;
    image[1][22][1] = 8'd144;
    image[1][22][2] = 8'd43;
    image[1][23][0] = 8'd49;
    image[1][23][1] = 8'd140;
    image[1][23][2] = 8'd40;
    image[1][24][0] = 8'd48;
    image[1][24][1] = 8'd138;
    image[1][24][2] = 8'd39;
    image[1][25][0] = 8'd49;
    image[1][25][1] = 8'd138;
    image[1][25][2] = 8'd39;
    image[1][26][0] = 8'd45;
    image[1][26][1] = 8'd133;
    image[1][26][2] = 8'd37;
    image[1][27][0] = 8'd45;
    image[1][27][1] = 8'd133;
    image[1][27][2] = 8'd37;
    image[1][28][0] = 8'd42;
    image[1][28][1] = 8'd130;
    image[1][28][2] = 8'd35;
    image[1][29][0] = 8'd41;
    image[1][29][1] = 8'd127;
    image[1][29][2] = 8'd35;
    image[2][0][0] = 8'd46;
    image[2][0][1] = 8'd131;
    image[2][0][2] = 8'd33;
    image[2][1][0] = 8'd45;
    image[2][1][1] = 8'd133;
    image[2][1][2] = 8'd34;
    image[2][2][0] = 8'd47;
    image[2][2][1] = 8'd135;
    image[2][2][2] = 8'd34;
    image[2][3][0] = 8'd47;
    image[2][3][1] = 8'd135;
    image[2][3][2] = 8'd35;
    image[2][4][0] = 8'd49;
    image[2][4][1] = 8'd138;
    image[2][4][2] = 8'd35;
    image[2][5][0] = 8'd49;
    image[2][5][1] = 8'd140;
    image[2][5][2] = 8'd34;
    image[2][6][0] = 8'd51;
    image[2][6][1] = 8'd143;
    image[2][6][2] = 8'd36;
    image[2][7][0] = 8'd51;
    image[2][7][1] = 8'd144;
    image[2][7][2] = 8'd36;
    image[2][8][0] = 8'd53;
    image[2][8][1] = 8'd146;
    image[2][8][2] = 8'd38;
    image[2][9][0] = 8'd54;
    image[2][9][1] = 8'd148;
    image[2][9][2] = 8'd38;
    image[2][10][0] = 8'd53;
    image[2][10][1] = 8'd149;
    image[2][10][2] = 8'd39;
    image[2][11][0] = 8'd52;
    image[2][11][1] = 8'd148;
    image[2][11][2] = 8'd37;
    image[2][12][0] = 8'd52;
    image[2][12][1] = 8'd148;
    image[2][12][2] = 8'd37;
    image[2][13][0] = 8'd55;
    image[2][13][1] = 8'd152;
    image[2][13][2] = 8'd41;
    image[2][14][0] = 8'd54;
    image[2][14][1] = 8'd150;
    image[2][14][2] = 8'd40;
    image[2][15][0] = 8'd51;
    image[2][15][1] = 8'd145;
    image[2][15][2] = 8'd38;
    image[2][16][0] = 8'd48;
    image[2][16][1] = 8'd140;
    image[2][16][2] = 8'd36;
    image[2][17][0] = 8'd48;
    image[2][17][1] = 8'd138;
    image[2][17][2] = 8'd36;
    image[2][18][0] = 8'd45;
    image[2][18][1] = 8'd136;
    image[2][18][2] = 8'd34;
    image[2][19][0] = 8'd47;
    image[2][19][1] = 8'd137;
    image[2][19][2] = 8'd37;
    image[2][20][0] = 8'd47;
    image[2][20][1] = 8'd136;
    image[2][20][2] = 8'd36;
    image[2][21][0] = 8'd49;
    image[2][21][1] = 8'd138;
    image[2][21][2] = 8'd37;
    image[2][22][0] = 8'd52;
    image[2][22][1] = 8'd141;
    image[2][22][2] = 8'd40;
    image[2][23][0] = 8'd52;
    image[2][23][1] = 8'd142;
    image[2][23][2] = 8'd41;
    image[2][24][0] = 8'd49;
    image[2][24][1] = 8'd140;
    image[2][24][2] = 8'd40;
    image[2][25][0] = 8'd47;
    image[2][25][1] = 8'd137;
    image[2][25][2] = 8'd38;
    image[2][26][0] = 8'd48;
    image[2][26][1] = 8'd137;
    image[2][26][2] = 8'd39;
    image[2][27][0] = 8'd46;
    image[2][27][1] = 8'd134;
    image[2][27][2] = 8'd37;
    image[2][28][0] = 8'd46;
    image[2][28][1] = 8'd133;
    image[2][28][2] = 8'd39;
    image[2][29][0] = 8'd42;
    image[2][29][1] = 8'd128;
    image[2][29][2] = 8'd36;
    image[3][0][0] = 8'd45;
    image[3][0][1] = 8'd133;
    image[3][0][2] = 8'd35;
    image[3][1][0] = 8'd45;
    image[3][1][1] = 8'd132;
    image[3][1][2] = 8'd33;
    image[3][2][0] = 8'd46;
    image[3][2][1] = 8'd135;
    image[3][2][2] = 8'd34;
    image[3][3][0] = 8'd50;
    image[3][3][1] = 8'd139;
    image[3][3][2] = 8'd36;
    image[3][4][0] = 8'd51;
    image[3][4][1] = 8'd140;
    image[3][4][2] = 8'd37;
    image[3][5][0] = 8'd53;
    image[3][5][1] = 8'd143;
    image[3][5][2] = 8'd38;
    image[3][6][0] = 8'd53;
    image[3][6][1] = 8'd144;
    image[3][6][2] = 8'd37;
    image[3][7][0] = 8'd53;
    image[3][7][1] = 8'd145;
    image[3][7][2] = 8'd37;
    image[3][8][0] = 8'd53;
    image[3][8][1] = 8'd148;
    image[3][8][2] = 8'd37;
    image[3][9][0] = 8'd53;
    image[3][9][1] = 8'd148;
    image[3][9][2] = 8'd37;
    image[3][10][0] = 8'd53;
    image[3][10][1] = 8'd150;
    image[3][10][2] = 8'd38;
    image[3][11][0] = 8'd55;
    image[3][11][1] = 8'd151;
    image[3][11][2] = 8'd39;
    image[3][12][0] = 8'd57;
    image[3][12][1] = 8'd153;
    image[3][12][2] = 8'd42;
    image[3][13][0] = 8'd56;
    image[3][13][1] = 8'd153;
    image[3][13][2] = 8'd42;
    image[3][14][0] = 8'd52;
    image[3][14][1] = 8'd144;
    image[3][14][2] = 8'd38;
    image[3][15][0] = 8'd41;
    image[3][15][1] = 8'd131;
    image[3][15][2] = 8'd32;
    image[3][16][0] = 8'd42;
    image[3][16][1] = 8'd129;
    image[3][16][2] = 8'd34;
    image[3][17][0] = 8'd43;
    image[3][17][1] = 8'd129;
    image[3][17][2] = 8'd35;
    image[3][18][0] = 8'd41;
    image[3][18][1] = 8'd126;
    image[3][18][2] = 8'd35;
    image[3][19][0] = 8'd41;
    image[3][19][1] = 8'd126;
    image[3][19][2] = 8'd35;
    image[3][20][0] = 8'd42;
    image[3][20][1] = 8'd127;
    image[3][20][2] = 8'd36;
    image[3][21][0] = 8'd41;
    image[3][21][1] = 8'd125;
    image[3][21][2] = 8'd34;
    image[3][22][0] = 8'd39;
    image[3][22][1] = 8'd122;
    image[3][22][2] = 8'd32;
    image[3][23][0] = 8'd44;
    image[3][23][1] = 8'd129;
    image[3][23][2] = 8'd36;
    image[3][24][0] = 8'd46;
    image[3][24][1] = 8'd133;
    image[3][24][2] = 8'd37;
    image[3][25][0] = 8'd44;
    image[3][25][1] = 8'd131;
    image[3][25][2] = 8'd35;
    image[3][26][0] = 8'd43;
    image[3][26][1] = 8'd129;
    image[3][26][2] = 8'd33;
    image[3][27][0] = 8'd40;
    image[3][27][1] = 8'd124;
    image[3][27][2] = 8'd31;
    image[3][28][0] = 8'd38;
    image[3][28][1] = 8'd121;
    image[3][28][2] = 8'd31;
    image[3][29][0] = 8'd35;
    image[3][29][1] = 8'd115;
    image[3][29][2] = 8'd29;
    image[4][0][0] = 8'd49;
    image[4][0][1] = 8'd135;
    image[4][0][2] = 8'd37;
    image[4][1][0] = 8'd49;
    image[4][1][1] = 8'd136;
    image[4][1][2] = 8'd36;
    image[4][2][0] = 8'd52;
    image[4][2][1] = 8'd140;
    image[4][2][2] = 8'd37;
    image[4][3][0] = 8'd53;
    image[4][3][1] = 8'd143;
    image[4][3][2] = 8'd38;
    image[4][4][0] = 8'd51;
    image[4][4][1] = 8'd143;
    image[4][4][2] = 8'd37;
    image[4][5][0] = 8'd53;
    image[4][5][1] = 8'd144;
    image[4][5][2] = 8'd36;
    image[4][6][0] = 8'd54;
    image[4][6][1] = 8'd145;
    image[4][6][2] = 8'd38;
    image[4][7][0] = 8'd55;
    image[4][7][1] = 8'd149;
    image[4][7][2] = 8'd38;
    image[4][8][0] = 8'd56;
    image[4][8][1] = 8'd150;
    image[4][8][2] = 8'd40;
    image[4][9][0] = 8'd54;
    image[4][9][1] = 8'd151;
    image[4][9][2] = 8'd38;
    image[4][10][0] = 8'd55;
    image[4][10][1] = 8'd152;
    image[4][10][2] = 8'd39;
    image[4][11][0] = 8'd54;
    image[4][11][1] = 8'd153;
    image[4][11][2] = 8'd39;
    image[4][12][0] = 8'd58;
    image[4][12][1] = 8'd154;
    image[4][12][2] = 8'd43;
    image[4][13][0] = 8'd48;
    image[4][13][1] = 8'd142;
    image[4][13][2] = 8'd35;
    image[4][14][0] = 8'd37;
    image[4][14][1] = 8'd123;
    image[4][14][2] = 8'd31;
    image[4][15][0] = 8'd36;
    image[4][15][1] = 8'd113;
    image[4][15][2] = 8'd37;
    image[4][16][0] = 8'd37;
    image[4][16][1] = 8'd107;
    image[4][16][2] = 8'd48;
    image[4][17][0] = 8'd37;
    image[4][17][1] = 8'd94;
    image[4][17][2] = 8'd63;
    image[4][18][0] = 8'd52;
    image[4][18][1] = 8'd105;
    image[4][18][2] = 8'd82;
    image[4][19][0] = 8'd60;
    image[4][19][1] = 8'd112;
    image[4][19][2] = 8'd92;
    image[4][20][0] = 8'd56;
    image[4][20][1] = 8'd108;
    image[4][20][2] = 8'd85;
    image[4][21][0] = 8'd33;
    image[4][21][1] = 8'd94;
    image[4][21][2] = 8'd50;
    image[4][22][0] = 8'd32;
    image[4][22][1] = 8'd104;
    image[4][22][2] = 8'd34;
    image[4][23][0] = 8'd34;
    image[4][23][1] = 8'd108;
    image[4][23][2] = 8'd33;
    image[4][24][0] = 8'd35;
    image[4][24][1] = 8'd113;
    image[4][24][2] = 8'd30;
    image[4][25][0] = 8'd35;
    image[4][25][1] = 8'd114;
    image[4][25][2] = 8'd31;
    image[4][26][0] = 8'd36;
    image[4][26][1] = 8'd114;
    image[4][26][2] = 8'd31;
    image[4][27][0] = 8'd35;
    image[4][27][1] = 8'd112;
    image[4][27][2] = 8'd30;
    image[4][28][0] = 8'd31;
    image[4][28][1] = 8'd107;
    image[4][28][2] = 8'd30;
    image[4][29][0] = 8'd29;
    image[4][29][1] = 8'd104;
    image[4][29][2] = 8'd29;
    image[5][0][0] = 8'd34;
    image[5][0][1] = 8'd117;
    image[5][0][2] = 8'd22;
    image[5][1][0] = 8'd48;
    image[5][1][1] = 8'd136;
    image[5][1][2] = 8'd33;
    image[5][2][0] = 8'd52;
    image[5][2][1] = 8'd141;
    image[5][2][2] = 8'd37;
    image[5][3][0] = 8'd52;
    image[5][3][1] = 8'd142;
    image[5][3][2] = 8'd37;
    image[5][4][0] = 8'd54;
    image[5][4][1] = 8'd145;
    image[5][4][2] = 8'd37;
    image[5][5][0] = 8'd53;
    image[5][5][1] = 8'd145;
    image[5][5][2] = 8'd37;
    image[5][6][0] = 8'd56;
    image[5][6][1] = 8'd149;
    image[5][6][2] = 8'd38;
    image[5][7][0] = 8'd57;
    image[5][7][1] = 8'd151;
    image[5][7][2] = 8'd41;
    image[5][8][0] = 8'd60;
    image[5][8][1] = 8'd154;
    image[5][8][2] = 8'd42;
    image[5][9][0] = 8'd57;
    image[5][9][1] = 8'd153;
    image[5][9][2] = 8'd39;
    image[5][10][0] = 8'd58;
    image[5][10][1] = 8'd155;
    image[5][10][2] = 8'd42;
    image[5][11][0] = 8'd59;
    image[5][11][1] = 8'd156;
    image[5][11][2] = 8'd43;
    image[5][12][0] = 8'd54;
    image[5][12][1] = 8'd149;
    image[5][12][2] = 8'd39;
    image[5][13][0] = 8'd42;
    image[5][13][1] = 8'd128;
    image[5][13][2] = 8'd34;
    image[5][14][0] = 8'd20;
    image[5][14][1] = 8'd85;
    image[5][14][2] = 8'd38;
    image[5][15][0] = 8'd97;
    image[5][15][1] = 8'd140;
    image[5][15][2] = 8'd153;
    image[5][16][0] = 8'd110;
    image[5][16][1] = 8'd144;
    image[5][16][2] = 8'd177;
    image[5][17][0] = 8'd88;
    image[5][17][1] = 8'd121;
    image[5][17][2] = 8'd157;
    image[5][18][0] = 8'd82;
    image[5][18][1] = 8'd116;
    image[5][18][2] = 8'd149;
    image[5][19][0] = 8'd77;
    image[5][19][1] = 8'd111;
    image[5][19][2] = 8'd143;
    image[5][20][0] = 8'd87;
    image[5][20][1] = 8'd119;
    image[5][20][2] = 8'd153;
    image[5][21][0] = 8'd87;
    image[5][21][1] = 8'd120;
    image[5][21][2] = 8'd152;
    image[5][22][0] = 8'd85;
    image[5][22][1] = 8'd120;
    image[5][22][2] = 8'd144;
    image[5][23][0] = 8'd66;
    image[5][23][1] = 8'd105;
    image[5][23][2] = 8'd113;
    image[5][24][0] = 8'd21;
    image[5][24][1] = 8'd75;
    image[5][24][2] = 8'd43;
    image[5][25][0] = 8'd15;
    image[5][25][1] = 8'd71;
    image[5][25][2] = 8'd33;
    image[5][26][0] = 8'd10;
    image[5][26][1] = 8'd65;
    image[5][26][2] = 8'd23;
    image[5][27][0] = 8'd12;
    image[5][27][1] = 8'd67;
    image[5][27][2] = 8'd24;
    image[5][28][0] = 8'd13;
    image[5][28][1] = 8'd67;
    image[5][28][2] = 8'd31;
    image[5][29][0] = 8'd15;
    image[5][29][1] = 8'd62;
    image[5][29][2] = 8'd33;
    image[6][0][0] = 8'd79;
    image[6][0][1] = 8'd158;
    image[6][0][2] = 8'd68;
    image[6][1][0] = 8'd57;
    image[6][1][1] = 8'd143;
    image[6][1][2] = 8'd42;
    image[6][2][0] = 8'd51;
    image[6][2][1] = 8'd142;
    image[6][2][2] = 8'd36;
    image[6][3][0] = 8'd54;
    image[6][3][1] = 8'd145;
    image[6][3][2] = 8'd37;
    image[6][4][0] = 8'd55;
    image[6][4][1] = 8'd146;
    image[6][4][2] = 8'd38;
    image[6][5][0] = 8'd55;
    image[6][5][1] = 8'd148;
    image[6][5][2] = 8'd38;
    image[6][6][0] = 8'd58;
    image[6][6][1] = 8'd152;
    image[6][6][2] = 8'd41;
    image[6][7][0] = 8'd57;
    image[6][7][1] = 8'd152;
    image[6][7][2] = 8'd40;
    image[6][8][0] = 8'd56;
    image[6][8][1] = 8'd153;
    image[6][8][2] = 8'd40;
    image[6][9][0] = 8'd58;
    image[6][9][1] = 8'd156;
    image[6][9][2] = 8'd40;
    image[6][10][0] = 8'd58;
    image[6][10][1] = 8'd156;
    image[6][10][2] = 8'd40;
    image[6][11][0] = 8'd58;
    image[6][11][1] = 8'd156;
    image[6][11][2] = 8'd42;
    image[6][12][0] = 8'd44;
    image[6][12][1] = 8'd138;
    image[6][12][2] = 8'd33;
    image[6][13][0] = 8'd36;
    image[6][13][1] = 8'd118;
    image[6][13][2] = 8'd34;
    image[6][14][0] = 8'd39;
    image[6][14][1] = 8'd91;
    image[6][14][2] = 8'd74;
    image[6][15][0] = 8'd122;
    image[6][15][1] = 8'd158;
    image[6][15][2] = 8'd189;
    image[6][16][0] = 8'd124;
    image[6][16][1] = 8'd155;
    image[6][16][2] = 8'd192;
    image[6][17][0] = 8'd109;
    image[6][17][1] = 8'd140;
    image[6][17][2] = 8'd179;
    image[6][18][0] = 8'd112;
    image[6][18][1] = 8'd143;
    image[6][18][2] = 8'd180;
    image[6][19][0] = 8'd105;
    image[6][19][1] = 8'd137;
    image[6][19][2] = 8'd175;
    image[6][20][0] = 8'd87;
    image[6][20][1] = 8'd120;
    image[6][20][2] = 8'd157;
    image[6][21][0] = 8'd100;
    image[6][21][1] = 8'd133;
    image[6][21][2] = 8'd169;
    image[6][22][0] = 8'd57;
    image[6][22][1] = 8'd91;
    image[6][22][2] = 8'd124;
    image[6][23][0] = 8'd70;
    image[6][23][1] = 8'd103;
    image[6][23][2] = 8'd134;
    image[6][24][0] = 8'd76;
    image[6][24][1] = 8'd110;
    image[6][24][2] = 8'd140;
    image[6][25][0] = 8'd90;
    image[6][25][1] = 8'd123;
    image[6][25][2] = 8'd155;
    image[6][26][0] = 8'd78;
    image[6][26][1] = 8'd110;
    image[6][26][2] = 8'd142;
    image[6][27][0] = 8'd91;
    image[6][27][1] = 8'd123;
    image[6][27][2] = 8'd158;
    image[6][28][0] = 8'd85;
    image[6][28][1] = 8'd118;
    image[6][28][2] = 8'd147;
    image[6][29][0] = 8'd63;
    image[6][29][1] = 8'd96;
    image[6][29][2] = 8'd121;
    image[7][0][0] = 8'd42;
    image[7][0][1] = 8'd127;
    image[7][0][2] = 8'd26;
    image[7][1][0] = 8'd54;
    image[7][1][1] = 8'd146;
    image[7][1][2] = 8'd37;
    image[7][2][0] = 8'd55;
    image[7][2][1] = 8'd148;
    image[7][2][2] = 8'd37;
    image[7][3][0] = 8'd54;
    image[7][3][1] = 8'd146;
    image[7][3][2] = 8'd37;
    image[7][4][0] = 8'd53;
    image[7][4][1] = 8'd146;
    image[7][4][2] = 8'd36;
    image[7][5][0] = 8'd54;
    image[7][5][1] = 8'd148;
    image[7][5][2] = 8'd36;
    image[7][6][0] = 8'd58;
    image[7][6][1] = 8'd152;
    image[7][6][2] = 8'd42;
    image[7][7][0] = 8'd56;
    image[7][7][1] = 8'd152;
    image[7][7][2] = 8'd39;
    image[7][8][0] = 8'd56;
    image[7][8][1] = 8'd153;
    image[7][8][2] = 8'd39;
    image[7][9][0] = 8'd56;
    image[7][9][1] = 8'd154;
    image[7][9][2] = 8'd39;
    image[7][10][0] = 8'd60;
    image[7][10][1] = 8'd158;
    image[7][10][2] = 8'd42;
    image[7][11][0] = 8'd55;
    image[7][11][1] = 8'd153;
    image[7][11][2] = 8'd40;
    image[7][12][0] = 8'd43;
    image[7][12][1] = 8'd133;
    image[7][12][2] = 8'd33;
    image[7][13][0] = 8'd27;
    image[7][13][1] = 8'd101;
    image[7][13][2] = 8'd35;
    image[7][14][0] = 8'd34;
    image[7][14][1] = 8'd81;
    image[7][14][2] = 8'd82;
    image[7][15][0] = 8'd108;
    image[7][15][1] = 8'd142;
    image[7][15][2] = 8'd181;
    image[7][16][0] = 8'd118;
    image[7][16][1] = 8'd150;
    image[7][16][2] = 8'd190;
    image[7][17][0] = 8'd122;
    image[7][17][1] = 8'd153;
    image[7][17][2] = 8'd192;
    image[7][18][0] = 8'd125;
    image[7][18][1] = 8'd157;
    image[7][18][2] = 8'd193;
    image[7][19][0] = 8'd126;
    image[7][19][1] = 8'd157;
    image[7][19][2] = 8'd193;
    image[7][20][0] = 8'd114;
    image[7][20][1] = 8'd147;
    image[7][20][2] = 8'd183;
    image[7][21][0] = 8'd84;
    image[7][21][1] = 8'd118;
    image[7][21][2] = 8'd154;
    image[7][22][0] = 8'd98;
    image[7][22][1] = 8'd131;
    image[7][22][2] = 8'd167;
    image[7][23][0] = 8'd95;
    image[7][23][1] = 8'd128;
    image[7][23][2] = 8'd164;
    image[7][24][0] = 8'd104;
    image[7][24][1] = 8'd137;
    image[7][24][2] = 8'd171;
    image[7][25][0] = 8'd104;
    image[7][25][1] = 8'd136;
    image[7][25][2] = 8'd171;
    image[7][26][0] = 8'd77;
    image[7][26][1] = 8'd108;
    image[7][26][2] = 8'd144;
    image[7][27][0] = 8'd92;
    image[7][27][1] = 8'd124;
    image[7][27][2] = 8'd160;
    image[7][28][0] = 8'd67;
    image[7][28][1] = 8'd99;
    image[7][28][2] = 8'd133;
    image[7][29][0] = 8'd95;
    image[7][29][1] = 8'd126;
    image[7][29][2] = 8'd160;
    image[8][0][0] = 8'd57;
    image[8][0][1] = 8'd143;
    image[8][0][2] = 8'd45;
    image[8][1][0] = 8'd55;
    image[8][1][1] = 8'd148;
    image[8][1][2] = 8'd39;
    image[8][2][0] = 8'd53;
    image[8][2][1] = 8'd147;
    image[8][2][2] = 8'd37;
    image[8][3][0] = 8'd54;
    image[8][3][1] = 8'd147;
    image[8][3][2] = 8'd37;
    image[8][4][0] = 8'd55;
    image[8][4][1] = 8'd148;
    image[8][4][2] = 8'd36;
    image[8][5][0] = 8'd55;
    image[8][5][1] = 8'd151;
    image[8][5][2] = 8'd38;
    image[8][6][0] = 8'd56;
    image[8][6][1] = 8'd152;
    image[8][6][2] = 8'd40;
    image[8][7][0] = 8'd58;
    image[8][7][1] = 8'd155;
    image[8][7][2] = 8'd41;
    image[8][8][0] = 8'd59;
    image[8][8][1] = 8'd156;
    image[8][8][2] = 8'd43;
    image[8][9][0] = 8'd57;
    image[8][9][1] = 8'd156;
    image[8][9][2] = 8'd40;
    image[8][10][0] = 8'd63;
    image[8][10][1] = 8'd161;
    image[8][10][2] = 8'd46;
    image[8][11][0] = 8'd52;
    image[8][11][1] = 8'd149;
    image[8][11][2] = 8'd39;
    image[8][12][0] = 8'd37;
    image[8][12][1] = 8'd122;
    image[8][12][2] = 8'd31;
    image[8][13][0] = 8'd25;
    image[8][13][1] = 8'd85;
    image[8][13][2] = 8'd47;
    image[8][14][0] = 8'd105;
    image[8][14][1] = 8'd145;
    image[8][14][2] = 8'd175;
    image[8][15][0] = 8'd147;
    image[8][15][1] = 8'd181;
    image[8][15][2] = 8'd217;
    image[8][16][0] = 8'd115;
    image[8][16][1] = 8'd147;
    image[8][16][2] = 8'd186;
    image[8][17][0] = 8'd111;
    image[8][17][1] = 8'd143;
    image[8][17][2] = 8'd180;
    image[8][18][0] = 8'd102;
    image[8][18][1] = 8'd134;
    image[8][18][2] = 8'd169;
    image[8][19][0] = 8'd115;
    image[8][19][1] = 8'd146;
    image[8][19][2] = 8'd180;
    image[8][20][0] = 8'd112;
    image[8][20][1] = 8'd144;
    image[8][20][2] = 8'd178;
    image[8][21][0] = 8'd106;
    image[8][21][1] = 8'd140;
    image[8][21][2] = 8'd175;
    image[8][22][0] = 8'd94;
    image[8][22][1] = 8'd128;
    image[8][22][2] = 8'd164;
    image[8][23][0] = 8'd102;
    image[8][23][1] = 8'd136;
    image[8][23][2] = 8'd174;
    image[8][24][0] = 8'd93;
    image[8][24][1] = 8'd129;
    image[8][24][2] = 8'd166;
    image[8][25][0] = 8'd88;
    image[8][25][1] = 8'd123;
    image[8][25][2] = 8'd161;
    image[8][26][0] = 8'd83;
    image[8][26][1] = 8'd119;
    image[8][26][2] = 8'd157;
    image[8][27][0] = 8'd85;
    image[8][27][1] = 8'd122;
    image[8][27][2] = 8'd159;
    image[8][28][0] = 8'd93;
    image[8][28][1] = 8'd129;
    image[8][28][2] = 8'd165;
    image[8][29][0] = 8'd77;
    image[8][29][1] = 8'd112;
    image[8][29][2] = 8'd149;
    image[9][0][0] = 8'd57;
    image[9][0][1] = 8'd142;
    image[9][0][2] = 8'd46;
    image[9][1][0] = 8'd53;
    image[9][1][1] = 8'd146;
    image[9][1][2] = 8'd37;
    image[9][2][0] = 8'd54;
    image[9][2][1] = 8'd147;
    image[9][2][2] = 8'd37;
    image[9][3][0] = 8'd54;
    image[9][3][1] = 8'd149;
    image[9][3][2] = 8'd38;
    image[9][4][0] = 8'd56;
    image[9][4][1] = 8'd151;
    image[9][4][2] = 8'd38;
    image[9][5][0] = 8'd55;
    image[9][5][1] = 8'd150;
    image[9][5][2] = 8'd37;
    image[9][6][0] = 8'd60;
    image[9][6][1] = 8'd155;
    image[9][6][2] = 8'd42;
    image[9][7][0] = 8'd58;
    image[9][7][1] = 8'd155;
    image[9][7][2] = 8'd42;
    image[9][8][0] = 8'd60;
    image[9][8][1] = 8'd157;
    image[9][8][2] = 8'd44;
    image[9][9][0] = 8'd61;
    image[9][9][1] = 8'd158;
    image[9][9][2] = 8'd45;
    image[9][10][0] = 8'd62;
    image[9][10][1] = 8'd159;
    image[9][10][2] = 8'd46;
    image[9][11][0] = 8'd43;
    image[9][11][1] = 8'd134;
    image[9][11][2] = 8'd32;
    image[9][12][0] = 8'd28;
    image[9][12][1] = 8'd104;
    image[9][12][2] = 8'd32;
    image[9][13][0] = 8'd44;
    image[9][13][1] = 8'd95;
    image[9][13][2] = 8'd85;
    image[9][14][0] = 8'd84;
    image[9][14][1] = 8'd126;
    image[9][14][2] = 8'd158;
    image[9][15][0] = 8'd108;
    image[9][15][1] = 8'd144;
    image[9][15][2] = 8'd181;
    image[9][16][0] = 8'd119;
    image[9][16][1] = 8'd151;
    image[9][16][2] = 8'd190;
    image[9][17][0] = 8'd109;
    image[9][17][1] = 8'd143;
    image[9][17][2] = 8'd178;
    image[9][18][0] = 8'd135;
    image[9][18][1] = 8'd167;
    image[9][18][2] = 8'd199;
    image[9][19][0] = 8'd135;
    image[9][19][1] = 8'd166;
    image[9][19][2] = 8'd197;
    image[9][20][0] = 8'd112;
    image[9][20][1] = 8'd144;
    image[9][20][2] = 8'd177;
    image[9][21][0] = 8'd125;
    image[9][21][1] = 8'd156;
    image[9][21][2] = 8'd189;
    image[9][22][0] = 8'd107;
    image[9][22][1] = 8'd139;
    image[9][22][2] = 8'd173;
    image[9][23][0] = 8'd89;
    image[9][23][1] = 8'd126;
    image[9][23][2] = 8'd163;
    image[9][24][0] = 8'd84;
    image[9][24][1] = 8'd121;
    image[9][24][2] = 8'd161;
    image[9][25][0] = 8'd101;
    image[9][25][1] = 8'd138;
    image[9][25][2] = 8'd176;
    image[9][26][0] = 8'd68;
    image[9][26][1] = 8'd104;
    image[9][26][2] = 8'd144;
    image[9][27][0] = 8'd74;
    image[9][27][1] = 8'd110;
    image[9][27][2] = 8'd149;
    image[9][28][0] = 8'd77;
    image[9][28][1] = 8'd113;
    image[9][28][2] = 8'd151;
    image[9][29][0] = 8'd84;
    image[9][29][1] = 8'd120;
    image[9][29][2] = 8'd158;
    image[10][0][0] = 8'd48;
    image[10][0][1] = 8'd131;
    image[10][0][2] = 8'd39;
    image[10][1][0] = 8'd53;
    image[10][1][1] = 8'd147;
    image[10][1][2] = 8'd36;
    image[10][2][0] = 8'd53;
    image[10][2][1] = 8'd147;
    image[10][2][2] = 8'd34;
    image[10][3][0] = 8'd56;
    image[10][3][1] = 8'd150;
    image[10][3][2] = 8'd39;
    image[10][4][0] = 8'd55;
    image[10][4][1] = 8'd150;
    image[10][4][2] = 8'd37;
    image[10][5][0] = 8'd56;
    image[10][5][1] = 8'd151;
    image[10][5][2] = 8'd38;
    image[10][6][0] = 8'd58;
    image[10][6][1] = 8'd154;
    image[10][6][2] = 8'd41;
    image[10][7][0] = 8'd56;
    image[10][7][1] = 8'd154;
    image[10][7][2] = 8'd40;
    image[10][8][0] = 8'd57;
    image[10][8][1] = 8'd155;
    image[10][8][2] = 8'd41;
    image[10][9][0] = 8'd60;
    image[10][9][1] = 8'd157;
    image[10][9][2] = 8'd43;
    image[10][10][0] = 8'd52;
    image[10][10][1] = 8'd147;
    image[10][10][2] = 8'd38;
    image[10][11][0] = 8'd40;
    image[10][11][1] = 8'd126;
    image[10][11][2] = 8'd36;
    image[10][12][0] = 8'd45;
    image[10][12][1] = 8'd104;
    image[10][12][2] = 8'd76;
    image[10][13][0] = 8'd53;
    image[10][13][1] = 8'd95;
    image[10][13][2] = 8'd113;
    image[10][14][0] = 8'd80;
    image[10][14][1] = 8'd118;
    image[10][14][2] = 8'd160;
    image[10][15][0] = 8'd158;
    image[10][15][1] = 8'd192;
    image[10][15][2] = 8'd230;
    image[10][16][0] = 8'd127;
    image[10][16][1] = 8'd162;
    image[10][16][2] = 8'd203;
    image[10][17][0] = 8'd134;
    image[10][17][1] = 8'd168;
    image[10][17][2] = 8'd204;
    image[10][18][0] = 8'd141;
    image[10][18][1] = 8'd175;
    image[10][18][2] = 8'd209;
    image[10][19][0] = 8'd138;
    image[10][19][1] = 8'd170;
    image[10][19][2] = 8'd205;
    image[10][20][0] = 8'd123;
    image[10][20][1] = 8'd157;
    image[10][20][2] = 8'd192;
    image[10][21][0] = 8'd121;
    image[10][21][1] = 8'd155;
    image[10][21][2] = 8'd189;
    image[10][22][0] = 8'd125;
    image[10][22][1] = 8'd161;
    image[10][22][2] = 8'd195;
    image[10][23][0] = 8'd106;
    image[10][23][1] = 8'd143;
    image[10][23][2] = 8'd179;
    image[10][24][0] = 8'd102;
    image[10][24][1] = 8'd141;
    image[10][24][2] = 8'd177;
    image[10][25][0] = 8'd105;
    image[10][25][1] = 8'd144;
    image[10][25][2] = 8'd180;
    image[10][26][0] = 8'd101;
    image[10][26][1] = 8'd139;
    image[10][26][2] = 8'd177;
    image[10][27][0] = 8'd80;
    image[10][27][1] = 8'd118;
    image[10][27][2] = 8'd157;
    image[10][28][0] = 8'd74;
    image[10][28][1] = 8'd111;
    image[10][28][2] = 8'd148;
    image[10][29][0] = 8'd67;
    image[10][29][1] = 8'd103;
    image[10][29][2] = 8'd141;
    image[11][0][0] = 8'd57;
    image[11][0][1] = 8'd142;
    image[11][0][2] = 8'd48;
    image[11][1][0] = 8'd52;
    image[11][1][1] = 8'd145;
    image[11][1][2] = 8'd35;
    image[11][2][0] = 8'd54;
    image[11][2][1] = 8'd149;
    image[11][2][2] = 8'd37;
    image[11][3][0] = 8'd55;
    image[11][3][1] = 8'd151;
    image[11][3][2] = 8'd38;
    image[11][4][0] = 8'd55;
    image[11][4][1] = 8'd149;
    image[11][4][2] = 8'd37;
    image[11][5][0] = 8'd54;
    image[11][5][1] = 8'd148;
    image[11][5][2] = 8'd36;
    image[11][6][0] = 8'd56;
    image[11][6][1] = 8'd154;
    image[11][6][2] = 8'd40;
    image[11][7][0] = 8'd57;
    image[11][7][1] = 8'd155;
    image[11][7][2] = 8'd41;
    image[11][8][0] = 8'd59;
    image[11][8][1] = 8'd157;
    image[11][8][2] = 8'd42;
    image[11][9][0] = 8'd60;
    image[11][9][1] = 8'd157;
    image[11][9][2] = 8'd44;
    image[11][10][0] = 8'd43;
    image[11][10][1] = 8'd138;
    image[11][10][2] = 8'd33;
    image[11][11][0] = 8'd38;
    image[11][11][1] = 8'd118;
    image[11][11][2] = 8'd40;
    image[11][12][0] = 8'd65;
    image[11][12][1] = 8'd108;
    image[11][12][2] = 8'd125;
    image[11][13][0] = 8'd52;
    image[11][13][1] = 8'd89;
    image[11][13][2] = 8'd120;
    image[11][14][0] = 8'd106;
    image[11][14][1] = 8'd144;
    image[11][14][2] = 8'd187;
    image[11][15][0] = 8'd141;
    image[11][15][1] = 8'd175;
    image[11][15][2] = 8'd212;
    image[11][16][0] = 8'd125;
    image[11][16][1] = 8'd158;
    image[11][16][2] = 8'd195;
    image[11][17][0] = 8'd139;
    image[11][17][1] = 8'd172;
    image[11][17][2] = 8'd207;
    image[11][18][0] = 8'd129;
    image[11][18][1] = 8'd162;
    image[11][18][2] = 8'd198;
    image[11][19][0] = 8'd106;
    image[11][19][1] = 8'd142;
    image[11][19][2] = 8'd178;
    image[11][20][0] = 8'd124;
    image[11][20][1] = 8'd159;
    image[11][20][2] = 8'd194;
    image[11][21][0] = 8'd134;
    image[11][21][1] = 8'd169;
    image[11][21][2] = 8'd205;
    image[11][22][0] = 8'd91;
    image[11][22][1] = 8'd127;
    image[11][22][2] = 8'd164;
    image[11][23][0] = 8'd92;
    image[11][23][1] = 8'd130;
    image[11][23][2] = 8'd170;
    image[11][24][0] = 8'd88;
    image[11][24][1] = 8'd127;
    image[11][24][2] = 8'd169;
    image[11][25][0] = 8'd87;
    image[11][25][1] = 8'd127;
    image[11][25][2] = 8'd169;
    image[11][26][0] = 8'd74;
    image[11][26][1] = 8'd112;
    image[11][26][2] = 8'd154;
    image[11][27][0] = 8'd70;
    image[11][27][1] = 8'd107;
    image[11][27][2] = 8'd147;
    image[11][28][0] = 8'd58;
    image[11][28][1] = 8'd92;
    image[11][28][2] = 8'd132;
    image[11][29][0] = 8'd68;
    image[11][29][1] = 8'd101;
    image[11][29][2] = 8'd140;
    image[12][0][0] = 8'd52;
    image[12][0][1] = 8'd135;
    image[12][0][2] = 8'd41;
    image[12][1][0] = 8'd53;
    image[12][1][1] = 8'd147;
    image[12][1][2] = 8'd36;
    image[12][2][0] = 8'd52;
    image[12][2][1] = 8'd147;
    image[12][2][2] = 8'd36;
    image[12][3][0] = 8'd53;
    image[12][3][1] = 8'd147;
    image[12][3][2] = 8'd36;
    image[12][4][0] = 8'd54;
    image[12][4][1] = 8'd148;
    image[12][4][2] = 8'd37;
    image[12][5][0] = 8'd55;
    image[12][5][1] = 8'd150;
    image[12][5][2] = 8'd37;
    image[12][6][0] = 8'd55;
    image[12][6][1] = 8'd151;
    image[12][6][2] = 8'd38;
    image[12][7][0] = 8'd56;
    image[12][7][1] = 8'd153;
    image[12][7][2] = 8'd40;
    image[12][8][0] = 8'd55;
    image[12][8][1] = 8'd152;
    image[12][8][2] = 8'd39;
    image[12][9][0] = 8'd58;
    image[12][9][1] = 8'd156;
    image[12][9][2] = 8'd43;
    image[12][10][0] = 8'd47;
    image[12][10][1] = 8'd139;
    image[12][10][2] = 8'd36;
    image[12][11][0] = 8'd20;
    image[12][11][1] = 8'd93;
    image[12][11][2] = 8'd29;
    image[12][12][0] = 8'd57;
    image[12][12][1] = 8'd98;
    image[12][12][2] = 8'd120;
    image[12][13][0] = 8'd48;
    image[12][13][1] = 8'd83;
    image[12][13][2] = 8'd118;
    image[12][14][0] = 8'd65;
    image[12][14][1] = 8'd99;
    image[12][14][2] = 8'd142;
    image[12][15][0] = 8'd139;
    image[12][15][1] = 8'd172;
    image[12][15][2] = 8'd206;
    image[12][16][0] = 8'd143;
    image[12][16][1] = 8'd175;
    image[12][16][2] = 8'd210;
    image[12][17][0] = 8'd141;
    image[12][17][1] = 8'd171;
    image[12][17][2] = 8'd204;
    image[12][18][0] = 8'd129;
    image[12][18][1] = 8'd162;
    image[12][18][2] = 8'd196;
    image[12][19][0] = 8'd137;
    image[12][19][1] = 8'd171;
    image[12][19][2] = 8'd206;
    image[12][20][0] = 8'd114;
    image[12][20][1] = 8'd151;
    image[12][20][2] = 8'd190;
    image[12][21][0] = 8'd94;
    image[12][21][1] = 8'd131;
    image[12][21][2] = 8'd170;
    image[12][22][0] = 8'd93;
    image[12][22][1] = 8'd131;
    image[12][22][2] = 8'd171;
    image[12][23][0] = 8'd94;
    image[12][23][1] = 8'd133;
    image[12][23][2] = 8'd175;
    image[12][24][0] = 8'd81;
    image[12][24][1] = 8'd122;
    image[12][24][2] = 8'd164;
    image[12][25][0] = 8'd94;
    image[12][25][1] = 8'd135;
    image[12][25][2] = 8'd176;
    image[12][26][0] = 8'd69;
    image[12][26][1] = 8'd109;
    image[12][26][2] = 8'd148;
    image[12][27][0] = 8'd64;
    image[12][27][1] = 8'd101;
    image[12][27][2] = 8'd138;
    image[12][28][0] = 8'd64;
    image[12][28][1] = 8'd102;
    image[12][28][2] = 8'd137;
    image[12][29][0] = 8'd58;
    image[12][29][1] = 8'd94;
    image[12][29][2] = 8'd126;
    image[13][0][0] = 8'd33;
    image[13][0][1] = 8'd120;
    image[13][0][2] = 8'd20;
    image[13][1][0] = 8'd56;
    image[13][1][1] = 8'd146;
    image[13][1][2] = 8'd38;
    image[13][2][0] = 8'd54;
    image[13][2][1] = 8'd146;
    image[13][2][2] = 8'd36;
    image[13][3][0] = 8'd54;
    image[13][3][1] = 8'd148;
    image[13][3][2] = 8'd37;
    image[13][4][0] = 8'd56;
    image[13][4][1] = 8'd148;
    image[13][4][2] = 8'd38;
    image[13][5][0] = 8'd56;
    image[13][5][1] = 8'd151;
    image[13][5][2] = 8'd39;
    image[13][6][0] = 8'd56;
    image[13][6][1] = 8'd152;
    image[13][6][2] = 8'd40;
    image[13][7][0] = 8'd58;
    image[13][7][1] = 8'd153;
    image[13][7][2] = 8'd40;
    image[13][8][0] = 8'd60;
    image[13][8][1] = 8'd156;
    image[13][8][2] = 8'd43;
    image[13][9][0] = 8'd55;
    image[13][9][1] = 8'd151;
    image[13][9][2] = 8'd39;
    image[13][10][0] = 8'd49;
    image[13][10][1] = 8'd135;
    image[13][10][2] = 8'd40;
    image[13][11][0] = 8'd58;
    image[13][11][1] = 8'd115;
    image[13][11][2] = 8'd95;
    image[13][12][0] = 8'd64;
    image[13][12][1] = 8'd104;
    image[13][12][2] = 8'd132;
    image[13][13][0] = 8'd60;
    image[13][13][1] = 8'd96;
    image[13][13][2] = 8'd133;
    image[13][14][0] = 8'd98;
    image[13][14][1] = 8'd136;
    image[13][14][2] = 8'd180;
    image[13][15][0] = 8'd151;
    image[13][15][1] = 8'd184;
    image[13][15][2] = 8'd220;
    image[13][16][0] = 8'd156;
    image[13][16][1] = 8'd190;
    image[13][16][2] = 8'd223;
    image[13][17][0] = 8'd135;
    image[13][17][1] = 8'd168;
    image[13][17][2] = 8'd204;
    image[13][18][0] = 8'd117;
    image[13][18][1] = 8'd153;
    image[13][18][2] = 8'd191;
    image[13][19][0] = 8'd104;
    image[13][19][1] = 8'd140;
    image[13][19][2] = 8'd181;
    image[13][20][0] = 8'd94;
    image[13][20][1] = 8'd132;
    image[13][20][2] = 8'd172;
    image[13][21][0] = 8'd102;
    image[13][21][1] = 8'd139;
    image[13][21][2] = 8'd179;
    image[13][22][0] = 8'd86;
    image[13][22][1] = 8'd124;
    image[13][22][2] = 8'd166;
    image[13][23][0] = 8'd82;
    image[13][23][1] = 8'd120;
    image[13][23][2] = 8'd162;
    image[13][24][0] = 8'd78;
    image[13][24][1] = 8'd118;
    image[13][24][2] = 8'd155;
    image[13][25][0] = 8'd15;
    image[13][25][1] = 8'd55;
    image[13][25][2] = 8'd65;
    image[13][26][0] = 8'd23;
    image[13][26][1] = 8'd65;
    image[13][26][2] = 8'd71;
    image[13][27][0] = 8'd6;
    image[13][27][1] = 8'd46;
    image[13][27][2] = 8'd44;
    image[13][28][0] = 8'd1;
    image[13][28][1] = 8'd37;
    image[13][28][2] = 8'd30;
    image[13][29][0] = 8'd0;
    image[13][29][1] = 8'd26;
    image[13][29][2] = 8'd18;
    image[14][0][0] = 8'd65;
    image[14][0][1] = 8'd145;
    image[14][0][2] = 8'd55;
    image[14][1][0] = 8'd32;
    image[14][1][1] = 8'd116;
    image[14][1][2] = 8'd16;
    image[14][2][0] = 8'd52;
    image[14][2][1] = 8'd143;
    image[14][2][2] = 8'd36;
    image[14][3][0] = 8'd53;
    image[14][3][1] = 8'd145;
    image[14][3][2] = 8'd36;
    image[14][4][0] = 8'd54;
    image[14][4][1] = 8'd147;
    image[14][4][2] = 8'd37;
    image[14][5][0] = 8'd54;
    image[14][5][1] = 8'd148;
    image[14][5][2] = 8'd37;
    image[14][6][0] = 8'd55;
    image[14][6][1] = 8'd149;
    image[14][6][2] = 8'd37;
    image[14][7][0] = 8'd59;
    image[14][7][1] = 8'd154;
    image[14][7][2] = 8'd41;
    image[14][8][0] = 8'd60;
    image[14][8][1] = 8'd155;
    image[14][8][2] = 8'd42;
    image[14][9][0] = 8'd54;
    image[14][9][1] = 8'd148;
    image[14][9][2] = 8'd40;
    image[14][10][0] = 8'd33;
    image[14][10][1] = 8'd112;
    image[14][10][2] = 8'd31;
    image[14][11][0] = 8'd36;
    image[14][11][1] = 8'd85;
    image[14][11][2] = 8'd75;
    image[14][12][0] = 8'd71;
    image[14][12][1] = 8'd109;
    image[14][12][2] = 8'd142;
    image[14][13][0] = 8'd69;
    image[14][13][1] = 8'd103;
    image[14][13][2] = 8'd145;
    image[14][14][0] = 8'd107;
    image[14][14][1] = 8'd144;
    image[14][14][2] = 8'd190;
    image[14][15][0] = 8'd165;
    image[14][15][1] = 8'd198;
    image[14][15][2] = 8'd234;
    image[14][16][0] = 8'd137;
    image[14][16][1] = 8'd171;
    image[14][16][2] = 8'd210;
    image[14][17][0] = 8'd101;
    image[14][17][1] = 8'd134;
    image[14][17][2] = 8'd176;
    image[14][18][0] = 8'd117;
    image[14][18][1] = 8'd152;
    image[14][18][2] = 8'd194;
    image[14][19][0] = 8'd98;
    image[14][19][1] = 8'd133;
    image[14][19][2] = 8'd173;
    image[14][20][0] = 8'd101;
    image[14][20][1] = 8'd138;
    image[14][20][2] = 8'd176;
    image[14][21][0] = 8'd104;
    image[14][21][1] = 8'd140;
    image[14][21][2] = 8'd177;
    image[14][22][0] = 8'd62;
    image[14][22][1] = 8'd101;
    image[14][22][2] = 8'd130;
    image[14][23][0] = 8'd36;
    image[14][23][1] = 8'd79;
    image[14][23][2] = 8'd90;
    image[14][24][0] = 8'd20;
    image[14][24][1] = 8'd81;
    image[14][24][2] = 8'd28;
    image[14][25][0] = 8'd28;
    image[14][25][1] = 8'd92;
    image[14][25][2] = 8'd29;
    image[14][26][0] = 8'd34;
    image[14][26][1] = 8'd103;
    image[14][26][2] = 8'd30;
    image[14][27][0] = 8'd34;
    image[14][27][1] = 8'd105;
    image[14][27][2] = 8'd28;
    image[14][28][0] = 8'd34;
    image[14][28][1] = 8'd106;
    image[14][28][2] = 8'd30;
    image[14][29][0] = 8'd28;
    image[14][29][1] = 8'd99;
    image[14][29][2] = 8'd26;
    image[15][0][0] = 8'd45;
    image[15][0][1] = 8'd131;
    image[15][0][2] = 8'd30;
    image[15][1][0] = 8'd51;
    image[15][1][1] = 8'd137;
    image[15][1][2] = 8'd34;
    image[15][2][0] = 8'd52;
    image[15][2][1] = 8'd143;
    image[15][2][2] = 8'd35;
    image[15][3][0] = 8'd51;
    image[15][3][1] = 8'd143;
    image[15][3][2] = 8'd35;
    image[15][4][0] = 8'd55;
    image[15][4][1] = 8'd146;
    image[15][4][2] = 8'd36;
    image[15][5][0] = 8'd55;
    image[15][5][1] = 8'd149;
    image[15][5][2] = 8'd38;
    image[15][6][0] = 8'd54;
    image[15][6][1] = 8'd148;
    image[15][6][2] = 8'd37;
    image[15][7][0] = 8'd56;
    image[15][7][1] = 8'd152;
    image[15][7][2] = 8'd41;
    image[15][8][0] = 8'd59;
    image[15][8][1] = 8'd154;
    image[15][8][2] = 8'd41;
    image[15][9][0] = 8'd47;
    image[15][9][1] = 8'd138;
    image[15][9][2] = 8'd35;
    image[15][10][0] = 8'd38;
    image[15][10][1] = 8'd116;
    image[15][10][2] = 8'd38;
    image[15][11][0] = 8'd78;
    image[15][11][1] = 8'd119;
    image[15][11][2] = 8'd131;
    image[15][12][0] = 8'd48;
    image[15][12][1] = 8'd82;
    image[15][12][2] = 8'd116;
    image[15][13][0] = 8'd45;
    image[15][13][1] = 8'd77;
    image[15][13][2] = 8'd119;
    image[15][14][0] = 8'd85;
    image[15][14][1] = 8'd122;
    image[15][14][2] = 8'd171;
    image[15][15][0] = 8'd106;
    image[15][15][1] = 8'd143;
    image[15][15][2] = 8'd186;
    image[15][16][0] = 8'd104;
    image[15][16][1] = 8'd139;
    image[15][16][2] = 8'd185;
    image[15][17][0] = 8'd93;
    image[15][17][1] = 8'd127;
    image[15][17][2] = 8'd171;
    image[15][18][0] = 8'd86;
    image[15][18][1] = 8'd121;
    image[15][18][2] = 8'd163;
    image[15][19][0] = 8'd98;
    image[15][19][1] = 8'd136;
    image[15][19][2] = 8'd177;
    image[15][20][0] = 8'd95;
    image[15][20][1] = 8'd132;
    image[15][20][2] = 8'd169;
    image[15][21][0] = 8'd47;
    image[15][21][1] = 8'd88;
    image[15][21][2] = 8'd103;
    image[15][22][0] = 8'd23;
    image[15][22][1] = 8'd72;
    image[15][22][2] = 8'd54;
    image[15][23][0] = 8'd32;
    image[15][23][1] = 8'd98;
    image[15][23][2] = 8'd36;
    image[15][24][0] = 8'd36;
    image[15][24][1] = 8'd110;
    image[15][24][2] = 8'd30;
    image[15][25][0] = 8'd44;
    image[15][25][1] = 8'd123;
    image[15][25][2] = 8'd32;
    image[15][26][0] = 8'd44;
    image[15][26][1] = 8'd125;
    image[15][26][2] = 8'd32;
    image[15][27][0] = 8'd41;
    image[15][27][1] = 8'd123;
    image[15][27][2] = 8'd31;
    image[15][28][0] = 8'd40;
    image[15][28][1] = 8'd122;
    image[15][28][2] = 8'd31;
    image[15][29][0] = 8'd40;
    image[15][29][1] = 8'd119;
    image[15][29][2] = 8'd32;
    image[16][0][0] = 8'd46;
    image[16][0][1] = 8'd133;
    image[16][0][2] = 8'd33;
    image[16][1][0] = 8'd50;
    image[16][1][1] = 8'd138;
    image[16][1][2] = 8'd35;
    image[16][2][0] = 8'd50;
    image[16][2][1] = 8'd140;
    image[16][2][2] = 8'd35;
    image[16][3][0] = 8'd52;
    image[16][3][1] = 8'd143;
    image[16][3][2] = 8'd36;
    image[16][4][0] = 8'd54;
    image[16][4][1] = 8'd145;
    image[16][4][2] = 8'd37;
    image[16][5][0] = 8'd52;
    image[16][5][1] = 8'd145;
    image[16][5][2] = 8'd35;
    image[16][6][0] = 8'd55;
    image[16][6][1] = 8'd148;
    image[16][6][2] = 8'd37;
    image[16][7][0] = 8'd56;
    image[16][7][1] = 8'd151;
    image[16][7][2] = 8'd41;
    image[16][8][0] = 8'd56;
    image[16][8][1] = 8'd150;
    image[16][8][2] = 8'd40;
    image[16][9][0] = 8'd51;
    image[16][9][1] = 8'd142;
    image[16][9][2] = 8'd38;
    image[16][10][0] = 8'd45;
    image[16][10][1] = 8'd127;
    image[16][10][2] = 8'd43;
    image[16][11][0] = 8'd48;
    image[16][11][1] = 8'd93;
    image[16][11][2] = 8'd92;
    image[16][12][0] = 8'd102;
    image[16][12][1] = 8'd134;
    image[16][12][2] = 8'd168;
    image[16][13][0] = 8'd118;
    image[16][13][1] = 8'd145;
    image[16][13][2] = 8'd187;
    image[16][14][0] = 8'd98;
    image[16][14][1] = 8'd126;
    image[16][14][2] = 8'd171;
    image[16][15][0] = 8'd93;
    image[16][15][1] = 8'd120;
    image[16][15][2] = 8'd162;
    image[16][16][0] = 8'd88;
    image[16][16][1] = 8'd116;
    image[16][16][2] = 8'd157;
    image[16][17][0] = 8'd82;
    image[16][17][1] = 8'd113;
    image[16][17][2] = 8'd148;
    image[16][18][0] = 8'd67;
    image[16][18][1] = 8'd103;
    image[16][18][2] = 8'd137;
    image[16][19][0] = 8'd54;
    image[16][19][1] = 8'd92;
    image[16][19][2] = 8'd115;
    image[16][20][0] = 8'd43;
    image[16][20][1] = 8'd88;
    image[16][20][2] = 8'd88;
    image[16][21][0] = 8'd30;
    image[16][21][1] = 8'd94;
    image[16][21][2] = 8'd39;
    image[16][22][0] = 8'd36;
    image[16][22][1] = 8'd106;
    image[16][22][2] = 8'd35;
    image[16][23][0] = 8'd46;
    image[16][23][1] = 8'd126;
    image[16][23][2] = 8'd35;
    image[16][24][0] = 8'd53;
    image[16][24][1] = 8'd140;
    image[16][24][2] = 8'd39;
    image[16][25][0] = 8'd53;
    image[16][25][1] = 8'd141;
    image[16][25][2] = 8'd38;
    image[16][26][0] = 8'd51;
    image[16][26][1] = 8'd139;
    image[16][26][2] = 8'd37;
    image[16][27][0] = 8'd50;
    image[16][27][1] = 8'd139;
    image[16][27][2] = 8'd38;
    image[16][28][0] = 8'd48;
    image[16][28][1] = 8'd135;
    image[16][28][2] = 8'd37;
    image[16][29][0] = 8'd49;
    image[16][29][1] = 8'd134;
    image[16][29][2] = 8'd39;
    image[17][0][0] = 8'd43;
    image[17][0][1] = 8'd132;
    image[17][0][2] = 8'd29;
    image[17][1][0] = 8'd48;
    image[17][1][1] = 8'd136;
    image[17][1][2] = 8'd33;
    image[17][2][0] = 8'd48;
    image[17][2][1] = 8'd137;
    image[17][2][2] = 8'd32;
    image[17][3][0] = 8'd50;
    image[17][3][1] = 8'd140;
    image[17][3][2] = 8'd35;
    image[17][4][0] = 8'd51;
    image[17][4][1] = 8'd141;
    image[17][4][2] = 8'd36;
    image[17][5][0] = 8'd50;
    image[17][5][1] = 8'd143;
    image[17][5][2] = 8'd34;
    image[17][6][0] = 8'd52;
    image[17][6][1] = 8'd145;
    image[17][6][2] = 8'd35;
    image[17][7][0] = 8'd55;
    image[17][7][1] = 8'd149;
    image[17][7][2] = 8'd38;
    image[17][8][0] = 8'd56;
    image[17][8][1] = 8'd150;
    image[17][8][2] = 8'd40;
    image[17][9][0] = 8'd55;
    image[17][9][1] = 8'd149;
    image[17][9][2] = 8'd40;
    image[17][10][0] = 8'd51;
    image[17][10][1] = 8'd141;
    image[17][10][2] = 8'd40;
    image[17][11][0] = 8'd33;
    image[17][11][1] = 8'd111;
    image[17][11][2] = 8'd32;
    image[17][12][0] = 8'd28;
    image[17][12][1] = 8'd99;
    image[17][12][2] = 8'd34;
    image[17][13][0] = 8'd90;
    image[17][13][1] = 8'd130;
    image[17][13][2] = 8'd150;
    image[17][14][0] = 8'd99;
    image[17][14][1] = 8'd134;
    image[17][14][2] = 8'd171;
    image[17][15][0] = 8'd97;
    image[17][15][1] = 8'd132;
    image[17][15][2] = 8'd170;
    image[17][16][0] = 8'd100;
    image[17][16][1] = 8'd136;
    image[17][16][2] = 8'd172;
    image[17][17][0] = 8'd81;
    image[17][17][1] = 8'd116;
    image[17][17][2] = 8'd149;
    image[17][18][0] = 8'd86;
    image[17][18][1] = 8'd124;
    image[17][18][2] = 8'd153;
    image[17][19][0] = 8'd37;
    image[17][19][1] = 8'd92;
    image[17][19][2] = 8'd62;
    image[17][20][0] = 8'd34;
    image[17][20][1] = 8'd106;
    image[17][20][2] = 8'd34;
    image[17][21][0] = 8'd42;
    image[17][21][1] = 8'd120;
    image[17][21][2] = 8'd34;
    image[17][22][0] = 8'd52;
    image[17][22][1] = 8'd137;
    image[17][22][2] = 8'd37;
    image[17][23][0] = 8'd54;
    image[17][23][1] = 8'd143;
    image[17][23][2] = 8'd40;
    image[17][24][0] = 8'd52;
    image[17][24][1] = 8'd141;
    image[17][24][2] = 8'd38;
    image[17][25][0] = 8'd52;
    image[17][25][1] = 8'd142;
    image[17][25][2] = 8'd39;
    image[17][26][0] = 8'd47;
    image[17][26][1] = 8'd138;
    image[17][26][2] = 8'd37;
    image[17][27][0] = 8'd50;
    image[17][27][1] = 8'd139;
    image[17][27][2] = 8'd39;
    image[17][28][0] = 8'd45;
    image[17][28][1] = 8'd134;
    image[17][28][2] = 8'd36;
    image[17][29][0] = 8'd45;
    image[17][29][1] = 8'd132;
    image[17][29][2] = 8'd37;
    image[18][0][0] = 8'd44;
    image[18][0][1] = 8'd131;
    image[18][0][2] = 8'd30;
    image[18][1][0] = 8'd46;
    image[18][1][1] = 8'd133;
    image[18][1][2] = 8'd31;
    image[18][2][0] = 8'd47;
    image[18][2][1] = 8'd136;
    image[18][2][2] = 8'd33;
    image[18][3][0] = 8'd47;
    image[18][3][1] = 8'd137;
    image[18][3][2] = 8'd32;
    image[18][4][0] = 8'd51;
    image[18][4][1] = 8'd141;
    image[18][4][2] = 8'd36;
    image[18][5][0] = 8'd49;
    image[18][5][1] = 8'd142;
    image[18][5][2] = 8'd34;
    image[18][6][0] = 8'd50;
    image[18][6][1] = 8'd143;
    image[18][6][2] = 8'd34;
    image[18][7][0] = 8'd55;
    image[18][7][1] = 8'd148;
    image[18][7][2] = 8'd38;
    image[18][8][0] = 8'd55;
    image[18][8][1] = 8'd149;
    image[18][8][2] = 8'd38;
    image[18][9][0] = 8'd55;
    image[18][9][1] = 8'd149;
    image[18][9][2] = 8'd37;
    image[18][10][0] = 8'd54;
    image[18][10][1] = 8'd149;
    image[18][10][2] = 8'd38;
    image[18][11][0] = 8'd54;
    image[18][11][1] = 8'd147;
    image[18][11][2] = 8'd40;
    image[18][12][0] = 8'd43;
    image[18][12][1] = 8'd129;
    image[18][12][2] = 8'd36;
    image[18][13][0] = 8'd39;
    image[18][13][1] = 8'd118;
    image[18][13][2] = 8'd38;
    image[18][14][0] = 8'd42;
    image[18][14][1] = 8'd119;
    image[18][14][2] = 8'd41;
    image[18][15][0] = 8'd37;
    image[18][15][1] = 8'd113;
    image[18][15][2] = 8'd34;
    image[18][16][0] = 8'd39;
    image[18][16][1] = 8'd116;
    image[18][16][2] = 8'd33;
    image[18][17][0] = 8'd43;
    image[18][17][1] = 8'd121;
    image[18][17][2] = 8'd36;
    image[18][18][0] = 8'd44;
    image[18][18][1] = 8'd123;
    image[18][18][2] = 8'd36;
    image[18][19][0] = 8'd44;
    image[18][19][1] = 8'd124;
    image[18][19][2] = 8'd35;
    image[18][20][0] = 8'd49;
    image[18][20][1] = 8'd133;
    image[18][20][2] = 8'd37;
    image[18][21][0] = 8'd53;
    image[18][21][1] = 8'd141;
    image[18][21][2] = 8'd38;
    image[18][22][0] = 8'd53;
    image[18][22][1] = 8'd145;
    image[18][22][2] = 8'd40;
    image[18][23][0] = 8'd51;
    image[18][23][1] = 8'd142;
    image[18][23][2] = 8'd37;
    image[18][24][0] = 8'd50;
    image[18][24][1] = 8'd141;
    image[18][24][2] = 8'd36;
    image[18][25][0] = 8'd50;
    image[18][25][1] = 8'd139;
    image[18][25][2] = 8'd36;
    image[18][26][0] = 8'd49;
    image[18][26][1] = 8'd137;
    image[18][26][2] = 8'd35;
    image[18][27][0] = 8'd47;
    image[18][27][1] = 8'd136;
    image[18][27][2] = 8'd36;
    image[18][28][0] = 8'd45;
    image[18][28][1] = 8'd133;
    image[18][28][2] = 8'd35;
    image[18][29][0] = 8'd44;
    image[18][29][1] = 8'd131;
    image[18][29][2] = 8'd36;
    image[19][0][0] = 8'd45;
    image[19][0][1] = 8'd130;
    image[19][0][2] = 8'd32;
    image[19][1][0] = 8'd45;
    image[19][1][1] = 8'd131;
    image[19][1][2] = 8'd31;
    image[19][2][0] = 8'd49;
    image[19][2][1] = 8'd136;
    image[19][2][2] = 8'd34;
    image[19][3][0] = 8'd48;
    image[19][3][1] = 8'd137;
    image[19][3][2] = 8'd32;
    image[19][4][0] = 8'd49;
    image[19][4][1] = 8'd139;
    image[19][4][2] = 8'd32;
    image[19][5][0] = 8'd49;
    image[19][5][1] = 8'd140;
    image[19][5][2] = 8'd33;
    image[19][6][0] = 8'd44;
    image[19][6][1] = 8'd137;
    image[19][6][2] = 8'd30;
    image[19][7][0] = 8'd50;
    image[19][7][1] = 8'd144;
    image[19][7][2] = 8'd35;
    image[19][8][0] = 8'd49;
    image[19][8][1] = 8'd145;
    image[19][8][2] = 8'd35;
    image[19][9][0] = 8'd49;
    image[19][9][1] = 8'd145;
    image[19][9][2] = 8'd34;
    image[19][10][0] = 8'd53;
    image[19][10][1] = 8'd149;
    image[19][10][2] = 8'd38;
    image[19][11][0] = 8'd53;
    image[19][11][1] = 8'd148;
    image[19][11][2] = 8'd37;
    image[19][12][0] = 8'd55;
    image[19][12][1] = 8'd149;
    image[19][12][2] = 8'd39;
    image[19][13][0] = 8'd52;
    image[19][13][1] = 8'd140;
    image[19][13][2] = 8'd39;
    image[19][14][0] = 8'd48;
    image[19][14][1] = 8'd135;
    image[19][14][2] = 8'd35;
    image[19][15][0] = 8'd51;
    image[19][15][1] = 8'd138;
    image[19][15][2] = 8'd38;
    image[19][16][0] = 8'd53;
    image[19][16][1] = 8'd140;
    image[19][16][2] = 8'd40;
    image[19][17][0] = 8'd53;
    image[19][17][1] = 8'd139;
    image[19][17][2] = 8'd38;
    image[19][18][0] = 8'd52;
    image[19][18][1] = 8'd138;
    image[19][18][2] = 8'd38;
    image[19][19][0] = 8'd55;
    image[19][19][1] = 8'd144;
    image[19][19][2] = 8'd39;
    image[19][20][0] = 8'd56;
    image[19][20][1] = 8'd145;
    image[19][20][2] = 8'd39;
    image[19][21][0] = 8'd52;
    image[19][21][1] = 8'd144;
    image[19][21][2] = 8'd36;
    image[19][22][0] = 8'd49;
    image[19][22][1] = 8'd142;
    image[19][22][2] = 8'd37;
    image[19][23][0] = 8'd51;
    image[19][23][1] = 8'd140;
    image[19][23][2] = 8'd36;
    image[19][24][0] = 8'd49;
    image[19][24][1] = 8'd139;
    image[19][24][2] = 8'd35;
    image[19][25][0] = 8'd47;
    image[19][25][1] = 8'd136;
    image[19][25][2] = 8'd33;
    image[19][26][0] = 8'd45;
    image[19][26][1] = 8'd133;
    image[19][26][2] = 8'd33;
    image[19][27][0] = 8'd46;
    image[19][27][1] = 8'd134;
    image[19][27][2] = 8'd34;
    image[19][28][0] = 8'd44;
    image[19][28][1] = 8'd132;
    image[19][28][2] = 8'd35;
    image[19][29][0] = 8'd43;
    image[19][29][1] = 8'd128;
    image[19][29][2] = 8'd34;
end
endmodule
