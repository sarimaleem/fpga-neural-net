`include "common.svh"

module data_init (input logic clk);

    logic [LENGTH-1][WIDTH-1] image;
    classifier classifier (clk, init_in, image);

    initial begin
        init_in = 0;
        image = 0;

        image[0][0] = 1'b0;
        image[0][1] = 1'b0;
        image[0][2] = 1'b0;
        image[0][3] = 1'b0;
        image[0][4] = 1'b0;
        image[0][5] = 1'b0;
        image[0][6] = 1'b0;
        image[0][7] = 1'b0;
        image[0][8] = 1'b0;
        image[0][9] = 1'b0;
        image[0][10] = 1'b0;
        image[0][11] = 1'b0;
        image[0][12] = 1'b0;
        image[0][13] = 1'b0;
        image[0][14] = 1'b0;
        image[0][15] = 1'b0;
        image[0][16] = 1'b0;
        image[0][17] = 1'b0;
        image[0][18] = 1'b0;
        image[0][19] = 1'b0;
        image[0][20] = 1'b0;
        image[0][21] = 1'b0;
        image[0][22] = 1'b0;
        image[0][23] = 1'b0;
        image[0][24] = 1'b0;
        image[0][25] = 1'b0;
        image[0][26] = 1'b0;
        image[0][27] = 1'b0;
        image[0][28] = 1'b0;
        image[0][29] = 1'b0;
        image[1][0] = 1'b0;
        image[1][1] = 1'b0;
        image[1][2] = 1'b0;
        image[1][3] = 1'b0;
        image[1][4] = 1'b0;
        image[1][5] = 1'b0;
        image[1][6] = 1'b0;
        image[1][7] = 1'b0;
        image[1][8] = 1'b0;
        image[1][9] = 1'b0;
        image[1][10] = 1'b0;
        image[1][11] = 1'b0;
        image[1][12] = 1'b0;
        image[1][13] = 1'b0;
        image[1][14] = 1'b0;
        image[1][15] = 1'b0;
        image[1][16] = 1'b0;
        image[1][17] = 1'b0;
        image[1][18] = 1'b0;
        image[1][19] = 1'b0;
        image[1][20] = 1'b0;
        image[1][21] = 1'b0;
        image[1][22] = 1'b0;
        image[1][23] = 1'b0;
        image[1][24] = 1'b0;
        image[1][25] = 1'b0;
        image[1][26] = 1'b0;
        image[1][27] = 1'b0;
        image[1][28] = 1'b0;
        image[1][29] = 1'b0;
        image[2][0] = 1'b0;
        image[2][1] = 1'b0;
        image[2][2] = 1'b0;
        image[2][3] = 1'b0;
        image[2][4] = 1'b0;
        image[2][5] = 1'b0;
        image[2][6] = 1'b0;
        image[2][7] = 1'b0;
        image[2][8] = 1'b0;
        image[2][9] = 1'b0;
        image[2][10] = 1'b0;
        image[2][11] = 1'b0;
        image[2][12] = 1'b0;
        image[2][13] = 1'b0;
        image[2][14] = 1'b0;
        image[2][15] = 1'b0;
        image[2][16] = 1'b0;
        image[2][17] = 1'b0;
        image[2][18] = 1'b0;
        image[2][19] = 1'b0;
        image[2][20] = 1'b0;
        image[2][21] = 1'b0;
        image[2][22] = 1'b0;
        image[2][23] = 1'b0;
        image[2][24] = 1'b0;
        image[2][25] = 1'b0;
        image[2][26] = 1'b0;
        image[2][27] = 1'b0;
        image[2][28] = 1'b0;
        image[2][29] = 1'b0;
        image[3][0] = 1'b0;
        image[3][1] = 1'b0;
        image[3][2] = 1'b0;
        image[3][3] = 1'b0;
        image[3][4] = 1'b0;
        image[3][5] = 1'b0;
        image[3][6] = 1'b0;
        image[3][7] = 1'b0;
        image[3][8] = 1'b0;
        image[3][9] = 1'b0;
        image[3][10] = 1'b0;
        image[3][11] = 1'b0;
        image[3][12] = 1'b0;
        image[3][13] = 1'b0;
        image[3][14] = 1'b0;
        image[3][15] = 1'b0;
        image[3][16] = 1'b0;
        image[3][17] = 1'b0;
        image[3][18] = 1'b0;
        image[3][19] = 1'b0;
        image[3][20] = 1'b0;
        image[3][21] = 1'b0;
        image[3][22] = 1'b0;
        image[3][23] = 1'b0;
        image[3][24] = 1'b0;
        image[3][25] = 1'b0;
        image[3][26] = 1'b0;
        image[3][27] = 1'b0;
        image[3][28] = 1'b0;
        image[3][29] = 1'b0;
        image[4][0] = 1'b0;
        image[4][1] = 1'b0;
        image[4][2] = 1'b0;
        image[4][3] = 1'b0;
        image[4][4] = 1'b0;
        image[4][5] = 1'b0;
        image[4][6] = 1'b0;
        image[4][7] = 1'b0;
        image[4][8] = 1'b0;
        image[4][9] = 1'b0;
        image[4][10] = 1'b0;
        image[4][11] = 1'b0;
        image[4][12] = 1'b0;
        image[4][13] = 1'b0;
        image[4][14] = 1'b0;
        image[4][15] = 1'b0;
        image[4][16] = 1'b0;
        image[4][17] = 1'b0;
        image[4][18] = 1'b0;
        image[4][19] = 1'b0;
        image[4][20] = 1'b0;
        image[4][21] = 1'b0;
        image[4][22] = 1'b0;
        image[4][23] = 1'b0;
        image[4][24] = 1'b0;
        image[4][25] = 1'b0;
        image[4][26] = 1'b0;
        image[4][27] = 1'b0;
        image[4][28] = 1'b0;
        image[4][29] = 1'b0;
        image[5][0] = 1'b0;
        image[5][1] = 1'b0;
        image[5][2] = 1'b0;
        image[5][3] = 1'b0;
        image[5][4] = 1'b0;
        image[5][5] = 1'b0;
        image[5][6] = 1'b0;
        image[5][7] = 1'b0;
        image[5][8] = 1'b0;
        image[5][9] = 1'b0;
        image[5][10] = 1'b0;
        image[5][11] = 1'b0;
        image[5][12] = 1'b0;
        image[5][13] = 1'b0;
        image[5][14] = 1'b0;
        image[5][15] = 1'b1;
        image[5][16] = 1'b1;
        image[5][17] = 1'b1;
        image[5][18] = 1'b1;
        image[5][19] = 1'b1;
        image[5][20] = 1'b1;
        image[5][21] = 1'b1;
        image[5][22] = 1'b1;
        image[5][23] = 1'b1;
        image[5][24] = 1'b0;
        image[5][25] = 1'b0;
        image[5][26] = 1'b0;
        image[5][27] = 1'b0;
        image[5][28] = 1'b0;
        image[5][29] = 1'b0;
        image[6][0] = 1'b0;
        image[6][1] = 1'b0;
        image[6][2] = 1'b0;
        image[6][3] = 1'b0;
        image[6][4] = 1'b0;
        image[6][5] = 1'b0;
        image[6][6] = 1'b0;
        image[6][7] = 1'b0;
        image[6][8] = 1'b0;
        image[6][9] = 1'b0;
        image[6][10] = 1'b0;
        image[6][11] = 1'b0;
        image[6][12] = 1'b0;
        image[6][13] = 1'b0;
        image[6][14] = 1'b0;
        image[6][15] = 1'b1;
        image[6][16] = 1'b1;
        image[6][17] = 1'b1;
        image[6][18] = 1'b1;
        image[6][19] = 1'b1;
        image[6][20] = 1'b1;
        image[6][21] = 1'b1;
        image[6][22] = 1'b1;
        image[6][23] = 1'b1;
        image[6][24] = 1'b1;
        image[6][25] = 1'b1;
        image[6][26] = 1'b1;
        image[6][27] = 1'b1;
        image[6][28] = 1'b1;
        image[6][29] = 1'b1;
        image[7][0] = 1'b0;
        image[7][1] = 1'b0;
        image[7][2] = 1'b0;
        image[7][3] = 1'b0;
        image[7][4] = 1'b0;
        image[7][5] = 1'b0;
        image[7][6] = 1'b0;
        image[7][7] = 1'b0;
        image[7][8] = 1'b0;
        image[7][9] = 1'b0;
        image[7][10] = 1'b0;
        image[7][11] = 1'b0;
        image[7][12] = 1'b0;
        image[7][13] = 1'b0;
        image[7][14] = 1'b1;
        image[7][15] = 1'b1;
        image[7][16] = 1'b1;
        image[7][17] = 1'b1;
        image[7][18] = 1'b1;
        image[7][19] = 1'b1;
        image[7][20] = 1'b1;
        image[7][21] = 1'b1;
        image[7][22] = 1'b1;
        image[7][23] = 1'b1;
        image[7][24] = 1'b1;
        image[7][25] = 1'b1;
        image[7][26] = 1'b1;
        image[7][27] = 1'b1;
        image[7][28] = 1'b1;
        image[7][29] = 1'b1;
        image[8][0] = 1'b0;
        image[8][1] = 1'b0;
        image[8][2] = 1'b0;
        image[8][3] = 1'b0;
        image[8][4] = 1'b0;
        image[8][5] = 1'b0;
        image[8][6] = 1'b0;
        image[8][7] = 1'b0;
        image[8][8] = 1'b0;
        image[8][9] = 1'b0;
        image[8][10] = 1'b0;
        image[8][11] = 1'b0;
        image[8][12] = 1'b0;
        image[8][13] = 1'b0;
        image[8][14] = 1'b1;
        image[8][15] = 1'b1;
        image[8][16] = 1'b1;
        image[8][17] = 1'b1;
        image[8][18] = 1'b1;
        image[8][19] = 1'b1;
        image[8][20] = 1'b1;
        image[8][21] = 1'b1;
        image[8][22] = 1'b1;
        image[8][23] = 1'b1;
        image[8][24] = 1'b1;
        image[8][25] = 1'b1;
        image[8][26] = 1'b1;
        image[8][27] = 1'b1;
        image[8][28] = 1'b1;
        image[8][29] = 1'b1;
        image[9][0] = 1'b0;
        image[9][1] = 1'b0;
        image[9][2] = 1'b0;
        image[9][3] = 1'b0;
        image[9][4] = 1'b0;
        image[9][5] = 1'b0;
        image[9][6] = 1'b0;
        image[9][7] = 1'b0;
        image[9][8] = 1'b0;
        image[9][9] = 1'b0;
        image[9][10] = 1'b0;
        image[9][11] = 1'b0;
        image[9][12] = 1'b0;
        image[9][13] = 1'b0;
        image[9][14] = 1'b1;
        image[9][15] = 1'b1;
        image[9][16] = 1'b1;
        image[9][17] = 1'b1;
        image[9][18] = 1'b1;
        image[9][19] = 1'b1;
        image[9][20] = 1'b1;
        image[9][21] = 1'b1;
        image[9][22] = 1'b1;
        image[9][23] = 1'b1;
        image[9][24] = 1'b1;
        image[9][25] = 1'b1;
        image[9][26] = 1'b1;
        image[9][27] = 1'b1;
        image[9][28] = 1'b1;
        image[9][29] = 1'b1;
        image[10][0] = 1'b0;
        image[10][1] = 1'b0;
        image[10][2] = 1'b0;
        image[10][3] = 1'b0;
        image[10][4] = 1'b0;
        image[10][5] = 1'b0;
        image[10][6] = 1'b0;
        image[10][7] = 1'b0;
        image[10][8] = 1'b0;
        image[10][9] = 1'b0;
        image[10][10] = 1'b0;
        image[10][11] = 1'b0;
        image[10][12] = 1'b0;
        image[10][13] = 1'b1;
        image[10][14] = 1'b1;
        image[10][15] = 1'b1;
        image[10][16] = 1'b1;
        image[10][17] = 1'b1;
        image[10][18] = 1'b1;
        image[10][19] = 1'b1;
        image[10][20] = 1'b1;
        image[10][21] = 1'b1;
        image[10][22] = 1'b1;
        image[10][23] = 1'b1;
        image[10][24] = 1'b1;
        image[10][25] = 1'b1;
        image[10][26] = 1'b1;
        image[10][27] = 1'b1;
        image[10][28] = 1'b1;
        image[10][29] = 1'b1;
        image[11][0] = 1'b0;
        image[11][1] = 1'b0;
        image[11][2] = 1'b0;
        image[11][3] = 1'b0;
        image[11][4] = 1'b0;
        image[11][5] = 1'b0;
        image[11][6] = 1'b0;
        image[11][7] = 1'b0;
        image[11][8] = 1'b0;
        image[11][9] = 1'b0;
        image[11][10] = 1'b0;
        image[11][11] = 1'b0;
        image[11][12] = 1'b1;
        image[11][13] = 1'b1;
        image[11][14] = 1'b1;
        image[11][15] = 1'b1;
        image[11][16] = 1'b1;
        image[11][17] = 1'b1;
        image[11][18] = 1'b1;
        image[11][19] = 1'b1;
        image[11][20] = 1'b1;
        image[11][21] = 1'b1;
        image[11][22] = 1'b1;
        image[11][23] = 1'b1;
        image[11][24] = 1'b1;
        image[11][25] = 1'b1;
        image[11][26] = 1'b1;
        image[11][27] = 1'b1;
        image[11][28] = 1'b1;
        image[11][29] = 1'b1;
        image[12][0] = 1'b0;
        image[12][1] = 1'b0;
        image[12][2] = 1'b0;
        image[12][3] = 1'b0;
        image[12][4] = 1'b0;
        image[12][5] = 1'b0;
        image[12][6] = 1'b0;
        image[12][7] = 1'b0;
        image[12][8] = 1'b0;
        image[12][9] = 1'b0;
        image[12][10] = 1'b0;
        image[12][11] = 1'b0;
        image[12][12] = 1'b1;
        image[12][13] = 1'b1;
        image[12][14] = 1'b1;
        image[12][15] = 1'b1;
        image[12][16] = 1'b1;
        image[12][17] = 1'b1;
        image[12][18] = 1'b1;
        image[12][19] = 1'b1;
        image[12][20] = 1'b1;
        image[12][21] = 1'b1;
        image[12][22] = 1'b1;
        image[12][23] = 1'b1;
        image[12][24] = 1'b1;
        image[12][25] = 1'b1;
        image[12][26] = 1'b1;
        image[12][27] = 1'b1;
        image[12][28] = 1'b1;
        image[12][29] = 1'b1;
        image[13][0] = 1'b0;
        image[13][1] = 1'b0;
        image[13][2] = 1'b0;
        image[13][3] = 1'b0;
        image[13][4] = 1'b0;
        image[13][5] = 1'b0;
        image[13][6] = 1'b0;
        image[13][7] = 1'b0;
        image[13][8] = 1'b0;
        image[13][9] = 1'b0;
        image[13][10] = 1'b0;
        image[13][11] = 1'b0;
        image[13][12] = 1'b1;
        image[13][13] = 1'b1;
        image[13][14] = 1'b1;
        image[13][15] = 1'b1;
        image[13][16] = 1'b1;
        image[13][17] = 1'b1;
        image[13][18] = 1'b1;
        image[13][19] = 1'b1;
        image[13][20] = 1'b1;
        image[13][21] = 1'b1;
        image[13][22] = 1'b1;
        image[13][23] = 1'b1;
        image[13][24] = 1'b1;
        image[13][25] = 1'b1;
        image[13][26] = 1'b0;
        image[13][27] = 1'b0;
        image[13][28] = 1'b0;
        image[13][29] = 1'b0;
        image[14][0] = 1'b0;
        image[14][1] = 1'b0;
        image[14][2] = 1'b0;
        image[14][3] = 1'b0;
        image[14][4] = 1'b0;
        image[14][5] = 1'b0;
        image[14][6] = 1'b0;
        image[14][7] = 1'b0;
        image[14][8] = 1'b0;
        image[14][9] = 1'b0;
        image[14][10] = 1'b0;
        image[14][11] = 1'b0;
        image[14][12] = 1'b1;
        image[14][13] = 1'b1;
        image[14][14] = 1'b1;
        image[14][15] = 1'b1;
        image[14][16] = 1'b1;
        image[14][17] = 1'b1;
        image[14][18] = 1'b1;
        image[14][19] = 1'b1;
        image[14][20] = 1'b1;
        image[14][21] = 1'b1;
        image[14][22] = 1'b1;
        image[14][23] = 1'b1;
        image[14][24] = 1'b0;
        image[14][25] = 1'b0;
        image[14][26] = 1'b0;
        image[14][27] = 1'b0;
        image[14][28] = 1'b0;
        image[14][29] = 1'b0;
        image[15][0] = 1'b0;
        image[15][1] = 1'b0;
        image[15][2] = 1'b0;
        image[15][3] = 1'b0;
        image[15][4] = 1'b0;
        image[15][5] = 1'b0;
        image[15][6] = 1'b0;
        image[15][7] = 1'b0;
        image[15][8] = 1'b0;
        image[15][9] = 1'b0;
        image[15][10] = 1'b0;
        image[15][11] = 1'b1;
        image[15][12] = 1'b1;
        image[15][13] = 1'b1;
        image[15][14] = 1'b1;
        image[15][15] = 1'b1;
        image[15][16] = 1'b1;
        image[15][17] = 1'b1;
        image[15][18] = 1'b1;
        image[15][19] = 1'b1;
        image[15][20] = 1'b1;
        image[15][21] = 1'b1;
        image[15][22] = 1'b0;
        image[15][23] = 1'b0;
        image[15][24] = 1'b0;
        image[15][25] = 1'b0;
        image[15][26] = 1'b0;
        image[15][27] = 1'b0;
        image[15][28] = 1'b0;
        image[15][29] = 1'b0;
        image[16][0] = 1'b0;
        image[16][1] = 1'b0;
        image[16][2] = 1'b0;
        image[16][3] = 1'b0;
        image[16][4] = 1'b0;
        image[16][5] = 1'b0;
        image[16][6] = 1'b0;
        image[16][7] = 1'b0;
        image[16][8] = 1'b0;
        image[16][9] = 1'b0;
        image[16][10] = 1'b0;
        image[16][11] = 1'b0;
        image[16][12] = 1'b1;
        image[16][13] = 1'b0;
        image[16][14] = 1'b0;
        image[16][15] = 1'b0;
        image[16][16] = 1'b0;
        image[16][17] = 1'b1;
        image[16][18] = 1'b1;
        image[16][19] = 1'b1;
        image[16][20] = 1'b0;
        image[16][21] = 1'b0;
        image[16][22] = 1'b0;
        image[16][23] = 1'b0;
        image[16][24] = 1'b0;
        image[16][25] = 1'b0;
        image[16][26] = 1'b0;
        image[16][27] = 1'b0;
        image[16][28] = 1'b0;
        image[16][29] = 1'b0;
        image[17][0] = 1'b0;
        image[17][1] = 1'b0;
        image[17][2] = 1'b0;
        image[17][3] = 1'b0;
        image[17][4] = 1'b0;
        image[17][5] = 1'b0;
        image[17][6] = 1'b0;
        image[17][7] = 1'b0;
        image[17][8] = 1'b0;
        image[17][9] = 1'b0;
        image[17][10] = 1'b0;
        image[17][11] = 1'b0;
        image[17][12] = 1'b0;
        image[17][13] = 1'b1;
        image[17][14] = 1'b1;
        image[17][15] = 1'b1;
        image[17][16] = 1'b1;
        image[17][17] = 1'b1;
        image[17][18] = 1'b1;
        image[17][19] = 1'b0;
        image[17][20] = 1'b0;
        image[17][21] = 1'b0;
        image[17][22] = 1'b0;
        image[17][23] = 1'b0;
        image[17][24] = 1'b0;
        image[17][25] = 1'b0;
        image[17][26] = 1'b0;
        image[17][27] = 1'b0;
        image[17][28] = 1'b0;
        image[17][29] = 1'b0;
        image[18][0] = 1'b0;
        image[18][1] = 1'b0;
        image[18][2] = 1'b0;
        image[18][3] = 1'b0;
        image[18][4] = 1'b0;
        image[18][5] = 1'b0;
        image[18][6] = 1'b0;
        image[18][7] = 1'b0;
        image[18][8] = 1'b0;
        image[18][9] = 1'b0;
        image[18][10] = 1'b0;
        image[18][11] = 1'b0;
        image[18][12] = 1'b0;
        image[18][13] = 1'b0;
        image[18][14] = 1'b0;
        image[18][15] = 1'b0;
        image[18][16] = 1'b0;
        image[18][17] = 1'b0;
        image[18][18] = 1'b0;
        image[18][19] = 1'b0;
        image[18][20] = 1'b0;
        image[18][21] = 1'b0;
        image[18][22] = 1'b0;
        image[18][23] = 1'b0;
        image[18][24] = 1'b0;
        image[18][25] = 1'b0;
        image[18][26] = 1'b0;
        image[18][27] = 1'b0;
        image[18][28] = 1'b0;
        image[18][29] = 1'b0;
        image[19][0] = 1'b0;
        image[19][1] = 1'b0;
        image[19][2] = 1'b0;
        image[19][3] = 1'b0;
        image[19][4] = 1'b0;
        image[19][5] = 1'b0;
        image[19][6] = 1'b0;
        image[19][7] = 1'b0;
        image[19][8] = 1'b0;
        image[19][9] = 1'b0;
        image[19][10] = 1'b0;
        image[19][11] = 1'b0;
        image[19][12] = 1'b0;
        image[19][13] = 1'b0;
        image[19][14] = 1'b0;
        image[19][15] = 1'b0;
        image[19][16] = 1'b0;
        image[19][17] = 1'b0;
        image[19][18] = 1'b0;
        image[19][19] = 1'b0;
        image[19][20] = 1'b0;
        image[19][21] = 1'b0;
        image[19][22] = 1'b0;
        image[19][23] = 1'b0;
        image[19][24] = 1'b0;
        image[19][25] = 1'b0;
        image[19][26] = 1'b0;
        image[19][27] = 1'b0;
        image[19][28] = 1'b0;
        image[19][29] = 1'b0;
    end
endmodule
